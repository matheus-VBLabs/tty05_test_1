

//IMPORTED BLOCK:bus_to_wires
// Bloco separador de barramento de 8 bits para uso na ferramenta 
module bus_to_wires (in,out_0,out_1,out_2,out_3,out_4,out_5,out_6,out_7);

// Inputs e Outputs
input wire [7:0] in;
output wire out_0,out_1,out_2,out_3,out_4,out_5,out_6,out_7;

// Comportamento do circuito
assign out_0 = in[0];
assign out_1 = in[1];
assign out_2 = in[2];
assign out_3 = in[3];
assign out_4 = in[4];
assign out_5 = in[5];
assign out_6 = in[6];
assign out_7 = in[7];

endmodule




//IMPORTED BLOCK:pulse_count_8_bits
module pulse_count_8_bits(pulse, counter);
input wire pulse;
output reg [7:0] counter;

initial counter = 0;

always @(posedge pulse) begin
counter <= counter + 1;
end

endmodule


// Automatically generated by ChipInventor Cloud EDA Tool - 2.0
// Careful: this file (hdl.v) will be automatically replaced when you ask
// to generate code from BLOCKS buttons.
module count_8_bits (

  input wire clk,
  output wire A3,
  output wire A4,
  output wire A2,
  output wire A5,
  output wire A1,
  output wire A6,
  output wire A8,
  output wire A7

);

//Internal Wires
 wire [7:0] w_1;

//Instances os Modules
pulse_count_8_bits blk82_20 (
         .pulse (clk),
         .counter (w_1)
     );

bus_to_wires blk28_22 (
         .out_2 (A3),
         .out_3 (A4),
         .out_1 (A2),
         .out_4 (A5),
         .out_0 (A1),
         .out_5 (A6),
         .out_7 (A8),
         .out_6 (A7),
         .in (w_1)
     );


endmodule
